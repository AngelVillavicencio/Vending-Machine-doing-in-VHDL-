library ieee;
use ieee.std_logic_1164.all;

entity bintobcd is
  port(signal a  :  in std_logic_vector(7 downto 0);
	   signal f  : out std_logic_vector(11 downto 0)) ;
end bintobcd;

architecture structural of bintobcd is

  constant DONT_CARE : std_logic_vector(11 downto 0):= (others => '-');

begin

  with a select
    f <= x"000" when x"00",
         x"001" when x"01",
         x"002" when x"02",
         x"003" when x"03",
         x"004" when x"04",
         x"005" when x"05",
         x"006" when x"06",
         x"007" when x"07",
         x"008" when x"08",
         x"009" when x"09",			 
         x"010" when x"0A",
         x"011" when x"0b",
         x"012" when x"0C",
         x"013" when x"0d",
         x"014" when x"0E",
         x"015" when x"0F",
         x"016" when x"10",
         x"017" when x"11",		 
         x"018" when x"12",
         x"019" when x"13",
         x"020" when x"14",	
         x"021" when x"15",
         x"022" when x"16",		 
         x"023" when x"17",
         x"024" when x"18",
         x"025" when x"19",	
         x"026" when x"1A",
         x"027" when x"1b",		 
         x"028" when x"1C",
         x"029" when x"1d",
         x"030" when x"1E",	
         x"031" when x"1F",	 
         x"032" when x"20",
         x"033" when x"21",
         x"034" when x"22",
         x"035" when x"23",
         x"036" when x"24",
         x"037" when x"25",
         x"038" when x"26",
         x"039" when x"27",
         x"040" when x"28",
         x"041" when x"29",			 
         x"042" when x"2A",
         x"043" when x"2b",
         x"044" when x"2C",
         x"045" when x"2d",
         x"046" when x"2E",
         x"047" when x"2F",
         x"048" when x"30",
         x"049" when x"31",		 
         x"050" when x"32",
         x"051" when x"33",
         x"052" when x"34",	
         x"053" when x"35",
         x"054" when x"36",		 
         x"055" when x"37",
         x"056" when x"38",
         x"057" when x"39",	
         x"058" when x"3A",
         x"059" when x"3b",		 
         x"060" when x"3C",
         x"061" when x"3D",
         x"062" when x"3E",	
         x"063" when x"3F",
         x"064" when x"40",
         x"065" when x"41",
         x"066" when x"42",
         x"067" when x"43",
         x"068" when x"44",
         x"069" when x"45",
         x"070" when x"46",
         x"071" when x"47",
         x"072" when x"48",
         x"073" when x"49",			 
         x"074" when x"4A",
         x"075" when x"4b",
         x"076" when x"4C",
         x"077" when x"4d",
         x"078" when x"4E",
         x"079" when x"4F",
         x"080" when x"50",
         x"081" when x"51",		 
         x"082" when x"52",
         x"083" when x"53",
         x"084" when x"54",	
         x"085" when x"55",
         x"086" when x"56",		 
         x"087" when x"57",
         x"088" when x"58",
         x"089" when x"59",	
         x"090" when x"5A",
         x"091" when x"5b",		 
         x"092" when x"5C",
         x"093" when x"5d",
         x"094" when x"5E",	
         x"095" when x"5F",
         x"096" when x"60",
         x"097" when x"61",
         x"098" when x"62",
         x"099" when x"63",
         x"100" when x"64",
         x"101" when x"65",
         x"102" when x"66",
         x"103" when x"67",
         x"104" when x"68",
         x"105" when x"69",			 
         x"106" when x"6A",
         x"107" when x"6b",
         x"108" when x"6C",
         x"109" when x"6d",
         x"110" when x"6E",
         x"111" when x"6F", 
         x"112" when x"70",
         x"113" when x"71",		 
         x"114" when x"72",
         x"115" when x"73",
         x"116" when x"74",	
         x"117" when x"75",
         x"118" when x"76",		 
         x"119" when x"77",
         x"120" when x"78",
         x"121" when x"79",	
         x"122" when x"7A",
         x"123" when x"7b",		 
         x"124" when x"7C",
         x"125" when x"7D",
         x"126" when x"7E",	
         x"127" when x"7F",		 
         x"128" when x"80",
         x"129" when x"81",		 
         x"130" when x"82",
         x"131" when x"83",
         x"132" when x"84",	
         x"133" when x"85",
         x"134" when x"86",		 
         x"135" when x"87",
         x"136" when x"88",
         x"137" when x"89",	
         x"138" when x"8A",
         x"139" when x"8b",		 
         x"140" when x"8C",
         x"141" when x"8D",
         x"142" when x"8E",	
         x"143" when x"8F",			 	 
         x"144" when x"90",
         x"145" when x"91",		 
         x"146" when x"92",
         x"147" when x"93",
         x"148" when x"94",	
         x"149" when x"95",
         x"150" when x"96",		 
         x"151" when x"97",
         x"152" when x"98",
         x"153" when x"99",	
         x"154" when x"9A",
         x"155" when x"9b",		 
         x"156" when x"9C",
         x"157" when x"9D",
         x"158" when x"9E",	
         x"159" when x"9F",		 	 
         x"160" when x"A0",
         x"161" when x"A1",		 
         x"162" when x"A2",
         x"163" when x"A3",
         x"164" when x"A4",	
         x"165" when x"A5",
         x"166" when x"A6",		 
         x"167" when x"A7",
         x"168" when x"A8",
         x"169" when x"A9",	
         x"170" when x"AA",
         x"171" when x"Ab",		 
         x"172" when x"AC",
         x"173" when x"AD",
         x"174" when x"AE",	
         x"175" when x"AF",		 
         x"176" when x"b0",
         x"177" when x"b1",		 
         x"178" when x"b2",
         x"179" when x"b3",
         x"180" when x"b4",	
         x"181" when x"b5",
         x"182" when x"b6",		 
         x"183" when x"b7",
         x"184" when x"b8",
         x"185" when x"b9",	
         x"186" when x"bA",
         x"187" when x"bb",		 
         x"188" when x"bC",
         x"189" when x"bD",
         x"190" when x"bE",	
         x"191" when x"bF",
         x"192" when x"C0",
         x"193" when x"C1",		 
         x"194" when x"C2",
         x"195" when x"C3",
         x"196" when x"C4",	
         x"197" when x"C5",
         x"198" when x"C6",		 
         x"199" when x"C7",
         x"200" when x"C8",
         x"201" when x"C9",	
         x"202" when x"CA",
         x"203" when x"Cb",		 
         x"204" when x"CC",
         x"205" when x"CD",
         x"206" when x"CE",	
         x"207" when x"CF",
         x"208" when x"D0",
         x"209" when x"D1",		 
         x"210" when x"D2",
         x"211" when x"D3",
         x"212" when x"D4",	
         x"213" when x"D5",
         x"214" when x"D6",		 
         x"215" when x"D7",
         x"216" when x"D8",
         x"217" when x"D9",	
         x"218" when x"DA",
         x"219" when x"Db",		 
         x"220" when x"DC",
         x"221" when x"DD",
         x"222" when x"DE",	
         x"223" when x"DF",
         x"224" when x"E0",
         x"225" when x"E1",		 
         x"226" when x"E2",
         x"227" when x"E3",
         x"228" when x"E4",	
         x"229" when x"E5",
         x"230" when x"E6",		 
         x"231" when x"E7",
         x"232" when x"E8",
         x"233" when x"E9",	
         x"234" when x"EA",
         x"235" when x"Eb",		 
         x"236" when x"EC",
         x"237" when x"ED",
         x"238" when x"EE",	
         x"239" when x"EF",
         x"240" when x"F0",
         x"241" when x"F1",		 
         x"242" when x"F2",
         x"243" when x"F3",
         x"244" when x"F4",	
         x"245" when x"F5",
         x"246" when x"F6",		 
         x"247" when x"F7",
         x"248" when x"F8",
         x"249" when x"F9",	
         x"250" when x"FA",
         x"251" when x"Fb",		 
         x"252" when x"FC",
         x"253" when x"FD",
         x"254" when x"FE",	
         x"255" when x"FF",
         DONT_CARE when others;

end structural;
